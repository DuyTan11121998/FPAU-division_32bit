module div_tb;
reg [31:0] A,B;

wire [31:0]S;

division uut(S,A,B);


initial begin
	A=32'h43d10000;
	B=32'h40000000;
#100
	A=32'h43800000;
	B=32'h42f00000;
#100
	A=32'h3f000000;
	B=32'h3e000000;
#100
	A=32'h3f000000;
	B=32'h41100000;
#100 
	A=32'h00000000;
	B=32'h00000000;
#100
	A=32'hc0c01100;
	B=32'h72800000;
#100
	A=32'hc0c00000;
	B=32'h74800000;
#100
	A=32'hc0c00000;
	B=32'h75800000;
#100
	A=32'hc0c00000;
	B=32'h1f800000;
#100
	A=32'hc0c00000;
	B=32'h4f800000;
#100
	A=32'hc0c00000;
	B=32'h5f800000;

end

endmodule
